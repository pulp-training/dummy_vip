`define DUMMY_SUCCESS_MESSAGE "Successfully integrated dummy IP."
